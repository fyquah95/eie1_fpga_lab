module adder(A,b,sum);
	input A[4:0];
	output B[4:0];
	
	assign sum = A + B;
	
endmodule